module glib

pub fn C.g_reload_user_special_dirs_cache()
pub fn g_reload_user_special_dirs_cache() {
	C.g_reload_user_special_dirs_cache()
}
