module glib

pub fn C.g_filesystem_preview_type_get_type() int
pub fn g_filesystem_preview_type_get_type() int {
	return C.g_filesystem_preview_type_get_type()
}
