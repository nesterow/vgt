module glib

pub fn C.g_password_save_get_type() int
pub fn g_password_save_get_type() int {
	return C.g_password_save_get_type()
}
