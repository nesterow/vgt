module glib

pub fn C.g_gtype_get_type() int
pub fn g_gtype_get_type() int {
	return C.g_gtype_get_type()
}
