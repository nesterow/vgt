module glib

pub fn C.g_blow_chunks()
pub fn g_blow_chunks() {
	C.g_blow_chunks()
}
