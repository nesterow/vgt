//
module main

import tool { GtkHeader, generate_gtk }

const frozen = true

fn main() {
	// 	// if frozen {
	// 	// 	println('codegen is frozen')
	// 	// 	return
	// 	// }

	// generate_gtk([GtkHeader{'gtkwidget', 'GtkWidget', 'gtk_widget', false}])!

	generate_gtk([
		GtkHeader{'gtkaboutdialog', 'GtkAboutDialog', 'gtk_about_dialog', false},
		GtkHeader{'gtkaccessible', 'GtkAccessible', 'gtk_accessible', false},
		GtkHeader{'gtkactionable', 'GtkActionable', 'gtk_actionable', false},
		GtkHeader{'gtkactionbar', 'GtkActionBar', 'gtk_action_bar', false},
		GtkHeader{'gtkadjustment', 'GtkAdjustment', 'gtk_adjustment', false},
		GtkHeader{'gtkappchooser', 'GtkAppChooser', 'gtk_app_chooser', false},
		GtkHeader{'gtkappchooserbutton', 'GtkAppChooserButton', 'gtk_app_chooser_button', false},
		GtkHeader{'gtkappchooserdialog', 'GtkAppChooserDialog', 'gtk_app_chooser_dialog', false},
		GtkHeader{'gtkappchooserwidget', 'GtkAppChooserWidget', 'gtk_app_chooser_widget', false},
		GtkHeader{'gtkapplication', 'GtkApplication', 'gtk_application', false},
		GtkHeader{'gtkapplicationwindow', 'GtkApplicationWindow', 'gtk_application_window', false},
		GtkHeader{'gtkaspectframe', 'GtkAspectFrame', 'gtk_aspect_frame', false},
		GtkHeader{'gtkassistant', 'GtkAssistant', 'gtk_assistant', false},
		GtkHeader{'gtkatcontext', 'GtkATContext', 'gtk_at_context', false},
		GtkHeader{'gtkbinlayout', 'GtkBinLayout', 'gtk_bin_layout', false},
		GtkHeader{'gtkbitset', 'GtkBitset', 'gtk_bitset', false},
		GtkHeader{'gtkbookmarklist', 'GtkBookmarkList', 'gtk_bookmark_list', false},
		GtkHeader{'gtkboolfilter', 'GtkBoolFilter', 'gtk_bool_filter', false},
		GtkHeader{'gtkborder', 'GtkBorder', 'gtk_border', false},
		GtkHeader{'gtkbox', 'GtkBox', 'gtk_box', false},
		GtkHeader{'gtkboxlayout', 'GtkBoxLayout', 'gtk_box_layout', false},
		GtkHeader{'gtkbuildable', 'GtkBuildable', 'gtk_buildable', false},
		GtkHeader{'gtkbuilder', 'GtkBuilderCScope', 'gtk_builder_cscope', false},
		GtkHeader{'gtkbuilder', 'GtkBuilder', 'gtk_builder', false},
		GtkHeader{'gtkbuilderlistitemfactory', 'GtkBuilderListItemFactory', 'gtk_builder_list_item_factory', false},
		GtkHeader{'gtkbutton', 'GtkButton', 'gtk_button', false},
		GtkHeader{'gtkcalendar', 'GtkCalendar', 'gtk_calendar', false},
		GtkHeader{'gtkcellarea', 'GtkCellArea', 'gtk_cell_area', false},
		GtkHeader{'gtkcellareabox', 'GtkCellAreaBox', 'gtk_cell_area_box', false},
		GtkHeader{'gtkcellareacontext', 'GtkCellAreaContext', 'gtk_cell_area_context', false},
		GtkHeader{'gtkcelleditable', 'GtkCellEditable', 'gtk_cell_editable', false},
		GtkHeader{'gtkcelllayout', 'GtkCellLayout', 'gtk_cell_layout', false},
		GtkHeader{'gtkcellrenderer', 'GtkCellRenderer', 'gtk_cell_renderer', false},
		GtkHeader{'gtkcellrendereraccel', 'GtkCellRendererAccel', 'gtk_cell_renderer_accel', false},
		GtkHeader{'gtkcellrenderercombo', 'GtkCellRendererCombo', 'gtk_cell_renderer_combo', false},
		GtkHeader{'gtkcellrendererpixbuf', 'GtkCellRendererPixbuf', 'gtk_cell_renderer_pixbuf', false},
		GtkHeader{'gtkcellrendererprogress', 'GtkCellRendererProgress', 'gtk_cell_renderer_progress', false},
		GtkHeader{'gtkcellrendererspin', 'GtkCellRendererSpin', 'gtk_cell_renderer_spin', false},
		GtkHeader{'gtkcellrendererspinner', 'GtkCellRendererSpinner', 'gtk_cell_renderer_spinner', false},
		GtkHeader{'gtkcellrenderertext', 'GtkCellRendererText', 'gtk_cell_renderer_text', false},
		GtkHeader{'gtkcellrenderertoggle', 'GtkCellRendererToggle', 'gtk_cell_renderer_toggle', false},
		GtkHeader{'gtkcellview', 'GtkCellView', 'gtk_cell_view', false},
		GtkHeader{'gtkcenterbox', 'GtkCenterBox', 'gtk_center_box', false},
		GtkHeader{'gtkcenterlayout', 'GtkCenterLayout', 'gtk_center_layout', false},
		GtkHeader{'gtkcheckbutton', 'GtkCheckButton', 'gtk_check_button', false},
		GtkHeader{'gtkcolorbutton', 'GtkColorButton', 'gtk_color_button', false},
		GtkHeader{'gtkcolorchooser', 'GtkColorChooser', 'gtk_color_chooser', false},
		GtkHeader{'gtkcolorchooserdialog', 'GtkColorChooserDialog', 'gtk_color_chooser_dialog', false},
		GtkHeader{'gtkcolorchooserwidget', 'GtkColorChooserWidget', 'gtk_color_chooser_widget', false},
		GtkHeader{'gtkcolumnview', 'GtkColumnView', 'gtk_column_view', false},
		GtkHeader{'gtkcolumnviewcolumn', 'GtkColumnViewColumn', 'gtk_column_view_column', false},
		GtkHeader{'gtkcombobox', 'GtkComboBox', 'gtk_combo_box', false},
		GtkHeader{'gtkcomboboxtext', 'GtkComboBoxText', 'gtk_combo_box_text', false},
		GtkHeader{'gtkconstraint', 'GtkConstraint', 'gtk_constraint', false},
		GtkHeader{'gtkconstraintguide', 'GtkConstraintGuide', 'gtk_constraint_guide', false},
		GtkHeader{'gtkconstraintlayout', 'GtkConstraintLayout', 'gtk_constraint_layout', false},
		GtkHeader{'gtkcssprovider', 'GtkCssProvider', 'gtk_css_provider', false},
		GtkHeader{'gtkcustomfilter', 'GtkCustomFilter', 'gtk_custom_filter', false},
		GtkHeader{'gtkcustomlayout', 'GtkCustomLayout', 'gtk_custom_layout', false},
		GtkHeader{'gtkcustomsorter', 'GtkCustomSorter', 'gtk_custom_sorter', false},
		GtkHeader{'gtkdialog', 'GtkDialog', 'gtk_dialog', false},
		GtkHeader{'gtkdirectorylist', 'GtkDirectoryList', 'gtk_directory_list', false},
		GtkHeader{'gtkdragicon', 'GtkDragIcon', 'gtk_drag_icon', false},
		GtkHeader{'gtkdragsource', 'GtkDragSource', 'gtk_drag_source', false},
		GtkHeader{'gtkdrawingarea', 'GtkDrawingArea', 'gtk_drawing_area', false},
		GtkHeader{'gtkdropcontrollermotion', 'GtkDropControllerMotion', 'gtk_drop_controller_motion', false},
		GtkHeader{'gtkdropdown', 'GtkDropDown', 'gtk_drop_down', false},
		GtkHeader{'gtkdroptarget', 'GtkDropTarget', 'gtk_drop_target', false},
		GtkHeader{'gtkdroptargetasync', 'GtkDropTargetAsync', 'gtk_drop_target_async', false},
		GtkHeader{'gtkeditable', 'GtkEditable', 'gtk_editable', false},
		GtkHeader{'gtkeditablelabel', 'GtkEditableLabel', 'gtk_editable_label', false},
		GtkHeader{'gtkemojichooser', 'GtkEmojiChooser', 'gtk_emoji_chooser', false},
		GtkHeader{'gtkentry', 'GtkEntry', 'gtk_entry', false},
		GtkHeader{'gtkentrybuffer', 'GtkEntryBuffer', 'gtk_entry_buffer', false},
		GtkHeader{'gtkentrycompletion', 'GtkEntryCompletion', 'gtk_entry_completion', false},
		GtkHeader{'gtkeventcontroller', 'GtkEventController', 'gtk_event_controller', false},
		GtkHeader{'gtkeventcontrollerfocus', 'GtkEventControllerFocus', 'gtk_event_controller_focus', false},
		GtkHeader{'gtkeventcontrollerkey', 'GtkEventControllerKey', 'gtk_event_controller_key', false},
		GtkHeader{'gtkeventcontrollermotion', 'GtkEventControllerMotion', 'gtk_event_controller_motion', false},
		GtkHeader{'gtkeventcontrollerscroll', 'GtkEventControllerScroll', 'gtk_event_controller_scroll', false},
		GtkHeader{'gtkexpander', 'GtkExpander', 'gtk_expander', false},
		GtkHeader{'gtkexpression', 'GtkExpression', 'gtk_expression', false},
		GtkHeader{'gtkfilechooser', 'GtkFileChooser', 'gtk_file_chooser', false},
		GtkHeader{'gtkfilechooserdialog', 'GtkFileChooserDialog', 'gtk_file_chooser_dialog', false},
		GtkHeader{'gtkfilechoosernative', 'GtkFileChooserNative', 'gtk_file_chooser_native', false},
		GtkHeader{'gtkfilechooserwidget', 'GtkFileChooserWidget', 'gtk_file_chooser_widget', false},
		GtkHeader{'gtkfilefilter', 'GtkFileFilter', 'gtk_file_filter', false},
		GtkHeader{'gtkfilter', 'GtkFilter', 'gtk_filter', false},
		GtkHeader{'gtkfilterlistmodel', 'GtkFilterListModel', 'gtk_filter_list_model', false},
		GtkHeader{'gtkfixed', 'GtkFixed', 'gtk_fixed', false},
		GtkHeader{'gtkfixedlayout', 'GtkFixedLayout', 'gtk_fixed_layout', false},
		GtkHeader{'gtkflattenlistmodel', 'GtkFlattenListModel', 'gtk_flatten_list_model', false},
		GtkHeader{'gtkflowbox', 'GtkFlowBoxChild', 'gtk_flow_box_child', false},
		GtkHeader{'gtkflowbox', 'GtkFlowBox', 'gtk_flow_box', false},
		GtkHeader{'gtkfontbutton', 'GtkFontButton', 'gtk_font_button', false},
		GtkHeader{'gtkfontchooser', 'GtkFontChooser', 'gtk_font_chooser', false},
		GtkHeader{'gtkfontchooserdialog', 'GtkFontChooserDialog', 'gtk_font_chooser_dialog', false},
		GtkHeader{'gtkfontchooserwidget', 'GtkFontChooserWidget', 'gtk_font_chooser_widget', false},
		GtkHeader{'gtkframe', 'GtkFrame', 'gtk_frame', false},
		GtkHeader{'gtkgesture', 'GtkGesture', 'gtk_gesture', false},
		GtkHeader{'gtkgestureclick', 'GtkGestureClick', 'gtk_gesture_click', false},
		GtkHeader{'gtkgesturedrag', 'GtkGestureDrag', 'gtk_gesture_drag', false},
		GtkHeader{'gtkgesturelongpress', 'GtkGestureLongPress', 'gtk_gesture_long_press', false},
		GtkHeader{'gtkgesturepan', 'GtkGesturePan', 'gtk_gesture_pan', false},
		GtkHeader{'gtkgesturerotate', 'GtkGestureRotate', 'gtk_gesture_rotate', false},
		GtkHeader{'gtkgesturesingle', 'GtkGestureSingle', 'gtk_gesture_single', false},
		GtkHeader{'gtkgesturestylus', 'GtkGestureStylus', 'gtk_gesture_stylus', false},
		GtkHeader{'gtkgestureswipe', 'GtkGestureSwipe', 'gtk_gesture_swipe', false},
		GtkHeader{'gtkgesturezoom', 'GtkGestureZoom', 'gtk_gesture_zoom', false},
		GtkHeader{'gtkglarea', 'GtkGLArea', 'gtk_gl_area', false},
		GtkHeader{'gtkgrid', 'GtkGrid', 'gtk_grid', false},
		GtkHeader{'gtkgridlayout', 'GtkGridLayout', 'gtk_grid_layout', false},
		GtkHeader{'gtkgridview', 'GtkGridView', 'gtk_grid_view', false},
		GtkHeader{'gtkheaderbar', 'GtkHeaderBar', 'gtk_header_bar', false},
		GtkHeader{'gtkicontheme', 'GtkIconPaintable', 'gtk_icon_paintable', false},
		GtkHeader{'gtkicontheme', 'GtkIconTheme', 'gtk_icon_theme', false},
		GtkHeader{'gtkiconview', 'GtkIconView', 'gtk_icon_view', false},
		GtkHeader{'gtkimage', 'GtkImage', 'gtk_image', false},
		GtkHeader{'gtkimcontext', 'GtkIMContext', 'gtk_im_context', false},
		GtkHeader{'gtkimcontextsimple', 'GtkIMContextSimple', 'gtk_im_context_simple', false},
		GtkHeader{'gtkimmulticontext', 'GtkIMMulticontext', 'gtk_im_multicontext', false},
		GtkHeader{'gtkinfobar', 'GtkInfoBar', 'gtk_info_bar', false},
		GtkHeader{'gtklabel', 'GtkLabel', 'gtk_label', false},
		GtkHeader{'gtklayoutchild', 'GtkLayoutChild', 'gtk_layout_child', false},
		GtkHeader{'gtklayoutmanager', 'GtkLayoutManager', 'gtk_layout_manager', false},
		GtkHeader{'gtklevelbar', 'GtkLevelBar', 'gtk_level_bar', false},
		GtkHeader{'gtklinkbutton', 'GtkLinkButton', 'gtk_link_button', false},
		GtkHeader{'gtklistbase', 'GtkListBase', 'gtk_list_base', false},
		GtkHeader{'gtklistbox', 'GtkListBox', 'gtk_list_box', false},
		GtkHeader{'gtklistitem', 'GtkListItem', 'gtk_list_item', false},
		GtkHeader{'gtklistitemfactory', 'GtkListItemFactory', 'gtk_list_item_factory', false},
		GtkHeader{'gtkliststore', 'GtkListStore', 'gtk_list_store', false},
		GtkHeader{'gtklistview', 'GtkListView', 'gtk_list_view', false},
		GtkHeader{'gtklockbutton', 'GtkLockButton', 'gtk_lock_button', false},
		GtkHeader{'gtkmaplistmodel', 'GtkMapListModel', 'gtk_map_list_model', false},
		GtkHeader{'gtkmediacontrols', 'GtkMediaControls', 'gtk_media_controls', false},
		GtkHeader{'gtkmediafile', 'GtkMediaFile', 'gtk_media_file', false},
		GtkHeader{'gtkmediastream', 'GtkMediaStream', 'gtk_media_stream', false},
		GtkHeader{'gtkmenubutton', 'GtkMenuButton', 'gtk_menu_button', false},
		GtkHeader{'gtkmessagedialog', 'GtkMessageDialog', 'gtk_message_dialog', false},
		GtkHeader{'gtkmountoperation', 'GtkMountOperation', 'gtk_mount_operation', false},
		GtkHeader{'gtkmultifilter', 'GtkMultiFilter', 'gtk_multi_filter', false},
		GtkHeader{'gtkmultiselection', 'GtkMultiSelection', 'gtk_multi_selection', false},
		GtkHeader{'gtkmultisorter', 'GtkMultiSorter', 'gtk_multi_sorter', false},
		GtkHeader{'gtknative', 'GtkNative', 'gtk_native', false},
		GtkHeader{'gtknativedialog', 'GtkNativeDialog', 'gtk_native_dialog', false},
		GtkHeader{'gtknoselection', 'GtkNoSelection', 'gtk_no_selection', false},
		GtkHeader{'gtknotebook', 'GtkNotebook', 'gtk_notebook', false},
		GtkHeader{'gtknumericsorter', 'GtkNumericSorter', 'gtk_numeric_sorter', false},
		GtkHeader{'gtkorientable', 'GtkOrientable', 'gtk_orientable', false},
		GtkHeader{'gtkoverlay', 'GtkOverlay', 'gtk_overlay', false},
		GtkHeader{'gtkoverlaylayout', 'GtkOverlayLayout', 'gtk_overlay_layout', false},
		GtkHeader{'gtkpadcontroller', 'GtkPadActionEntry', '$$', false},
		GtkHeader{'gtkpadcontroller', 'GtkPadController', 'gtk_pad_controller', false},
		GtkHeader{'gtkpagesetup', 'GtkPageSetup', 'gtk_page_setup', false},
		GtkHeader{'gtkpaned', 'GtkPaned', 'gtk_paned', false},
		GtkHeader{'gtkpapersize', 'GtkPaperSize', 'gtk_paper_size', false},
		GtkHeader{'gtkpasswordentry', 'GtkPasswordEntry', 'gtk_password_entry', false},
		GtkHeader{'gtkpasswordentrybuffer', 'GtkPasswordEntryBuffer', 'gtk_password_entry_buffer', false},
		GtkHeader{'gtkpicture', 'GtkPicture', 'gtk_picture', false},
		GtkHeader{'gtkpopover', 'GtkPopover', 'gtk_popover', false},
		GtkHeader{'gtkpopovermenu', 'GtkPopoverMenu', 'gtk_popover_menu', false},
		GtkHeader{'gtkpopovermenubar', 'GtkPopoverMenuBar', 'gtk_popover_menu_bar', false},
		GtkHeader{'gtkprintcontext', 'GtkPrintContext', 'gtk_print_context', false},
		GtkHeader{'gtkprintoperation', 'GtkPrintOperation', 'gtk_print_operation', false},
		GtkHeader{'gtkprintoperationpreview', 'GtkPrintOperationPreview', 'gtk_print_operation_preview', false},
		GtkHeader{'gtkprintsettings', 'GtkPrintSettings', 'gtk_print_settings', false},
		GtkHeader{'gtkprogressbar', 'GtkProgressBar', 'gtk_progress_bar', false},
		GtkHeader{'gtkrange', 'GtkRange', 'gtk_range', false},
		GtkHeader{'gtkrecentmanager', 'GtkRecentData', '$', false},
		GtkHeader{'gtkrecentmanager', 'GtkRecentInfo', '$', false},
		GtkHeader{'gtkrecentmanager', 'GtkRecentManager', 'gtk_recent_manager', false},
		GtkHeader{'gtkrevealer', 'GtkRevealer', 'gtk_revealer', false},
		GtkHeader{'gtkroot', 'GtkRoot', 'gtk_root', false},
		GtkHeader{'gtkscale', 'GtkScale', 'gtk_scale', false},
		GtkHeader{'gtkscalebutton', 'GtkScaleButton', 'gtk_scale_button', false},
		GtkHeader{'gtkscrollable', 'GtkScrollable', 'gtk_scrollable', false},
		GtkHeader{'gtkscrollbar', 'GtkScrollbar', 'gtk_scrollbar', false},
		GtkHeader{'gtkscrolledwindow', 'GtkScrolledWindow', 'gtk_scrolled_window', false},
		GtkHeader{'gtksearchbar', 'GtkSearchBar', 'gtk_search_bar', false},
		GtkHeader{'gtksearchentry', 'GtkSearchEntry', 'gtk_search_entry', false},
		GtkHeader{'gtkselectionfiltermodel', 'GtkSelectionModel', 'gtk_selection_model', false},
		GtkHeader{'gtkseparator', 'GtkSeparator', 'gtk_separator', false},
		GtkHeader{'gtksettings', 'GtkSettings', 'gtk_settings', false},
		GtkHeader{'gtkshortcut', 'GtkShortcut', 'gtk_shortcut', false},
		GtkHeader{'gtkshortcutaction', 'GtkShortcutAction', 'gtk_shortcut_action', false},
		GtkHeader{'gtkshortcutcontroller', 'GtkShortcutController', 'gtk_shortcut_controller', false},
		GtkHeader{'gtkshortcutlabel', 'GtkShortcutLabel', 'gtk_shortcut_label', false},
		GtkHeader{'gtkshortcutmanager', 'GtkShortcutManager', 'gtk_shortcut_manager', false},
		GtkHeader{'gtkshortcutsgroup', 'GtkShortcutsGroup', 'gtk_shortcuts_group', false},
		GtkHeader{'gtkshortcutssection', 'GtkShortcutsSection', 'gtk_shortcuts_section', false},
		GtkHeader{'gtkshortcutsshortcut', 'GtkShortcutsShortcut', 'gtk_shortcuts_shortcut', false},
		GtkHeader{'gtkshortcutswindow', 'GtkShortcutsWindow', 'gtk_shortcuts_window', false},
		GtkHeader{'gtkshortcuttrigger', 'GtkShortcutTrigger', 'gtk_shortcut_trigger', false},
		GtkHeader{'gtksignallistitemfactory', 'GtkSignalListItemFactory', 'gtk_signal_list_item_factory', false},
		GtkHeader{'gtksingleselection', 'GtkSingleSelection', 'gtk_single_selection', false},
		GtkHeader{'gtksizegroup', 'GtkSizeGroup', 'gtk_size_group', false},
		GtkHeader{'gtksizerequest', 'GtkRequestedSize', '$', false},
		GtkHeader{'gtkslicelistmodel', 'GtkSliceListModel', 'gtk_slice_list_model', false},
		GtkHeader{'gtksnapshot', 'GtkSnapshot', 'gtk_snapshot', false},
		GtkHeader{'gtksorter', 'GtkSorter', 'gtk_sorter', false},
		GtkHeader{'gtksortlistmodel', 'GtkSortListModel', 'gtk_sort_list_model', false},
		GtkHeader{'gtkspinbutton', 'GtkSpinButton', 'gtk_spin_button', false},
		GtkHeader{'gtkspinner', 'GtkSpinner', 'gtk_spinner', false},
		GtkHeader{'gtkstack', 'GtkStackPage', 'gtk_stack_page', false},
		GtkHeader{'gtkstack', 'GtkStack', 'gtk_stack', false},
		GtkHeader{'gtkstacksidebar', 'GtkStackSidebar', 'gtk_stack_sidebar', false},
		GtkHeader{'gtkstackswitcher', 'GtkStackSwitcher', 'gtk_stack_switcher', false},
		GtkHeader{'gtkstatusbar', 'GtkStatusbar', 'gtk_statusbar', false},
		GtkHeader{'gtkstringfilter', 'GtkStringFilter', 'gtk_string_filter', false},
		GtkHeader{'gtkstringlist', 'GtkStringList', 'gtk_string_list', false},
		GtkHeader{'gtkstringsorter', 'GtkStringSorter', 'gtk_string_sorter', false},
		GtkHeader{'gtkstylecontext', 'GtkStyleContext', 'gtk_style_context', false},
		GtkHeader{'gtkstyleprovider', 'GtkStyleProvider', 'gtk_style_provider', false},
		GtkHeader{'gtkswitch', 'GtkSwitch', 'gtk_switch', false},
		GtkHeader{'gtksymbolicpaintable', 'GtkSymbolicPaintable', 'gtk_symbolic_paintable', false},
		GtkHeader{'gtktext', 'GtkText', 'gtk_text', false},
		GtkHeader{'gtktextbuffer', 'GtkTextBuffer', 'gtk_text_buffer', false},
		GtkHeader{'gtktextchild', 'GtkTextChildAnchor', 'gtk_text_child', false},
		GtkHeader{'gtktextiter', 'GtkTextIter', 'gtk_text_iter', false},
		GtkHeader{'gtktextmark', 'GtkTextMark', 'gtk_text_mark', false},
		GtkHeader{'gtktexttag', 'GtkTextTag', 'gtk_text_tag', false},
		GtkHeader{'gtktexttagtable', 'GtkTextTagTable', 'gtk_text_tag_table', false},
		GtkHeader{'gtktextview', 'GtkTextView', 'gtk_text_view', false},
		GtkHeader{'gtktogglebutton', 'GtkToggleButton', 'gtk_toggle_button', false},
		GtkHeader{'gtktooltip', 'GtkTooltip', 'gtk_tooltip', false},
		GtkHeader{'gtktreednd', 'GtkTreeDragSource', 'gtk_tree_drag_source', false},
		GtkHeader{'gtktreednd', 'GtkTreeDragDest', 'gtk_tree_drag_dest', false},
		GtkHeader{'gtktreeexpander', 'GtkTreeExpander', 'gtk_tree_expander', false},
		GtkHeader{'gtktreelistmodel', 'GtkTreeListModel', 'gtk_tree_list_model', false},
		GtkHeader{'gtktreelistmodel', 'GtkTreeListRow', 'gtk_tree_list_row', false},
		GtkHeader{'gtktreelistrowsorter', 'GtkTreeListRowSorter', 'gtk_tree_list_row_sorter', false},
		GtkHeader{'gtktreemodel', 'GtkTreeModel', 'gtk_tree_model', false},
		GtkHeader{'gtktreemodel', 'GtkTreeIter', 'gtk_tree_iter', false},
		GtkHeader{'gtktreemodel', 'GtkTreePath', 'gtk_tree_path', false},
		GtkHeader{'gtktreemodel', 'GtkTreeRowReference', 'gtk_tree_row_reference', false},
		GtkHeader{'gtktreemodelfilter', 'GtkTreeModelFilter', 'gtk_tree_model_filter', false},
		GtkHeader{'gtktreemodelsort', 'GtkTreeModelSort', 'gtk_tree_model_sort', false},
		GtkHeader{'gtktreeselection', 'GtkTreeSelection', 'gtk_tree_selection', false},
		GtkHeader{'gtktreesortable', 'GtkTreeSortable', 'gtk_tree_sortable', false},
		GtkHeader{'gtktreestore', 'GtkTreeStore', 'gtk_tree_store', false},
		GtkHeader{'gtktreeviewcolumn', 'GtkTreeViewColumn', 'gtk_tree_view_column', false},
		GtkHeader{'gtktreeview', 'GtkTreeView', 'gtk_tree_view', false},
		GtkHeader{'gtkvideo', 'GtkVideo', 'gtk_video', false},
		GtkHeader{'gtkviewport', 'GtkViewport', 'gtk_viewport', false},
		GtkHeader{'gtkvolumebutton', 'GtkVolumeButton', 'gtk_volume_button', false},
		GtkHeader{'gtkwidget', 'GtkWidget', 'gtk_widget', false},
		GtkHeader{'gtkwindow', 'GtkWindow', 'gtk_window', false},
		GtkHeader{'gtkwidgetpaintable', 'GtkWidgetPaintable', 'gtk_widget_paintable', false},
		GtkHeader{'gtkwindowcontrols', 'GtkWindowControls', 'gtk_window_controls', false},
		GtkHeader{'gtkwindowgroup', 'GtkWindowGroup', 'gtk_window_group', false},
		GtkHeader{'gtkwindowhandle', 'GtkWindowHandle', 'gtk_window_handle', false},
	])!
}
