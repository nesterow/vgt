module glib

pub fn C.g_number_parser_error_quark() GQuark
pub fn g_number_parser_error_quark() GQuark {
	return C.g_number_parser_error_quark()
}
