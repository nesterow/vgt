module glib

pub fn C.g_normalize_mode_get_type() int
pub fn g_normalize_mode_get_type() int {
	return C.g_normalize_mode_get_type()
}
