module glib

pub fn C.g_ask_password_flags_get_type() int
pub fn g_ask_password_flags_get_type() int {
	return C.g_ask_password_flags_get_type()
}
