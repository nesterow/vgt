module glib

pub fn C.g_gstring_get_type() int
pub fn g_gstring_get_type() int {
	return C.g_gstring_get_type()
}
