module gtk
