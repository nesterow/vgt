module glib

pub fn C.g_unix_socket_address_type_get_type() int
pub fn g_unix_socket_address_type_get_type() int {
	return C.g_unix_socket_address_type_get_type()
}
