module glib

pub fn C.g_initially_unowned_get_type() int
pub fn g_initially_unowned_get_type() int {
	return C.g_initially_unowned_get_type()
}
