module gtk

@[noinit; typedef]
pub struct C.GtkRequestedSize {}

pub type GtkRequestedSize = C.GtkRequestedSize
